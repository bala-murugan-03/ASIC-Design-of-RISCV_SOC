VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbytes_1rw1r_20x256_20
   CLASS BLOCK ;
   SIZE 398.02 BY 392.565 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  76.54 0.0 76.92 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  82.38 0.0 82.76 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  88.22 0.0 88.6 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  94.06 0.0 94.44 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  99.9 0.0 100.28 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.74 0.0 106.12 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  111.58 0.0 111.96 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  117.42 0.0 117.8 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  123.26 0.0 123.64 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  129.1 0.0 129.48 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  134.94 0.0 135.32 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  140.78 0.0 141.16 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.62 0.0 147.0 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  152.46 0.0 152.84 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  158.3 0.0 158.68 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  164.14 0.0 164.52 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  169.98 0.0 170.36 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  175.82 0.0 176.2 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  181.66 0.0 182.04 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  187.5 0.0 187.88 0.38 ;
      END
   END din0[19]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.7 0.0 71.08 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 122.665 0.38 123.045 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 131.165 0.38 131.545 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.805 0.38 137.185 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 145.305 0.38 145.685 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 150.945 0.38 151.325 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 159.445 0.38 159.825 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 165.085 0.38 165.465 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  321.94 392.185 322.32 392.565 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.64 77.525 398.02 77.905 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.64 69.075 398.02 69.455 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.64 63.385 398.02 63.765 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  341.0 0.0 341.38 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  338.025 0.0 338.405 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  338.715 0.0 339.095 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  339.46 0.0 339.84 0.38 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 21.785 0.38 22.165 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  397.64 377.315 398.02 377.695 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 30.285 0.38 30.665 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  367.38 392.185 367.76 392.565 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  137.205 0.0 137.585 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.445 0.0 143.825 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  149.685 0.0 150.065 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.925 0.0 156.305 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.165 0.0 162.545 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  168.175 0.0 168.555 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.96 0.0 174.34 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  179.855 0.0 180.235 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  188.505 0.0 188.885 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.365 0.0 193.745 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.605 0.0 199.985 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.845 0.0 206.225 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.085 0.0 212.465 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.325 0.0 218.705 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.565 0.0 224.945 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.805 0.0 231.185 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  237.045 0.0 237.425 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  243.285 0.0 243.665 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  249.525 0.0 249.905 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.765 0.0 256.145 0.38 ;
      END
   END dout0[19]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  137.265 392.185 137.645 392.565 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.505 392.185 143.885 392.565 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  149.745 392.185 150.125 392.565 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.985 392.185 156.365 392.565 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.225 392.185 162.605 392.565 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  168.465 392.185 168.845 392.565 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  174.705 392.185 175.085 392.565 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.945 392.185 181.325 392.565 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.185 392.185 187.565 392.565 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.425 392.185 193.805 392.565 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  199.665 392.185 200.045 392.565 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  205.905 392.185 206.285 392.565 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.145 392.185 212.525 392.565 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.385 392.185 218.765 392.565 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.625 392.185 225.005 392.565 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.865 392.185 231.245 392.565 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  237.105 392.185 237.485 392.565 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  243.345 392.185 243.725 392.565 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  249.585 392.185 249.965 392.565 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  255.825 392.185 256.205 392.565 ;
      END
   END dout1[19]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 398.02 1.74 ;
         LAYER met3 ;
         RECT  0.0 390.825 398.02 392.565 ;
         LAYER met4 ;
         RECT  396.28 0.0 398.02 392.565 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 392.565 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.48 387.345 394.54 389.085 ;
         LAYER met3 ;
         RECT  3.48 3.48 394.54 5.22 ;
         LAYER met4 ;
         RECT  392.8 3.48 394.54 389.085 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 389.085 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 397.4 391.945 ;
   LAYER  met2 ;
      RECT  0.62 0.62 397.4 391.945 ;
   LAYER  met3 ;
      RECT  0.98 122.065 397.4 123.645 ;
      RECT  0.62 123.645 0.98 130.565 ;
      RECT  0.62 132.145 0.98 136.205 ;
      RECT  0.62 137.785 0.98 144.705 ;
      RECT  0.62 146.285 0.98 150.345 ;
      RECT  0.62 151.925 0.98 158.845 ;
      RECT  0.62 160.425 0.98 164.485 ;
      RECT  0.98 76.925 397.04 78.505 ;
      RECT  0.98 78.505 397.04 122.065 ;
      RECT  397.04 78.505 397.4 122.065 ;
      RECT  397.04 70.055 397.4 76.925 ;
      RECT  397.04 64.365 397.4 68.475 ;
      RECT  0.98 123.645 397.04 376.715 ;
      RECT  0.98 376.715 397.04 378.295 ;
      RECT  397.04 123.645 397.4 376.715 ;
      RECT  0.62 22.765 0.98 29.685 ;
      RECT  0.62 31.265 0.98 122.065 ;
      RECT  397.04 2.34 397.4 62.785 ;
      RECT  0.62 2.34 0.98 21.185 ;
      RECT  0.62 166.065 0.98 390.225 ;
      RECT  397.04 378.295 397.4 390.225 ;
      RECT  0.98 378.295 2.88 386.745 ;
      RECT  0.98 386.745 2.88 389.685 ;
      RECT  0.98 389.685 2.88 390.225 ;
      RECT  2.88 378.295 395.14 386.745 ;
      RECT  2.88 389.685 395.14 390.225 ;
      RECT  395.14 378.295 397.04 386.745 ;
      RECT  395.14 386.745 397.04 389.685 ;
      RECT  395.14 389.685 397.04 390.225 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 76.925 ;
      RECT  2.88 2.34 395.14 2.88 ;
      RECT  2.88 5.82 395.14 76.925 ;
      RECT  395.14 2.34 397.04 2.88 ;
      RECT  395.14 2.88 397.04 5.82 ;
      RECT  395.14 5.82 397.04 76.925 ;
   LAYER  met4 ;
      RECT  75.94 0.98 77.52 391.945 ;
      RECT  77.52 0.62 81.78 0.98 ;
      RECT  83.36 0.62 87.62 0.98 ;
      RECT  89.2 0.62 93.46 0.98 ;
      RECT  95.04 0.62 99.3 0.98 ;
      RECT  100.88 0.62 105.14 0.98 ;
      RECT  106.72 0.62 110.98 0.98 ;
      RECT  112.56 0.62 116.82 0.98 ;
      RECT  118.4 0.62 122.66 0.98 ;
      RECT  124.24 0.62 128.5 0.98 ;
      RECT  130.08 0.62 134.34 0.98 ;
      RECT  182.64 0.62 186.9 0.98 ;
      RECT  71.68 0.62 75.94 0.98 ;
      RECT  77.52 0.98 321.34 391.585 ;
      RECT  321.34 0.98 322.92 391.585 ;
      RECT  32.08 0.62 70.1 0.98 ;
      RECT  322.92 391.585 366.78 391.945 ;
      RECT  135.92 0.62 136.605 0.98 ;
      RECT  138.185 0.62 140.18 0.98 ;
      RECT  141.76 0.62 142.845 0.98 ;
      RECT  144.425 0.62 146.02 0.98 ;
      RECT  147.6 0.62 149.085 0.98 ;
      RECT  150.665 0.62 151.86 0.98 ;
      RECT  153.44 0.62 155.325 0.98 ;
      RECT  156.905 0.62 157.7 0.98 ;
      RECT  159.28 0.62 161.565 0.98 ;
      RECT  163.145 0.62 163.54 0.98 ;
      RECT  165.12 0.62 167.575 0.98 ;
      RECT  169.155 0.62 169.38 0.98 ;
      RECT  170.96 0.62 173.36 0.98 ;
      RECT  174.94 0.62 175.22 0.98 ;
      RECT  176.8 0.62 179.255 0.98 ;
      RECT  180.835 0.62 181.06 0.98 ;
      RECT  189.485 0.62 192.765 0.98 ;
      RECT  194.345 0.62 199.005 0.98 ;
      RECT  200.585 0.62 205.245 0.98 ;
      RECT  206.825 0.62 211.485 0.98 ;
      RECT  213.065 0.62 217.725 0.98 ;
      RECT  219.305 0.62 223.965 0.98 ;
      RECT  225.545 0.62 230.205 0.98 ;
      RECT  231.785 0.62 236.445 0.98 ;
      RECT  238.025 0.62 242.685 0.98 ;
      RECT  244.265 0.62 248.925 0.98 ;
      RECT  250.505 0.62 255.165 0.98 ;
      RECT  256.745 0.62 337.425 0.98 ;
      RECT  77.52 391.585 136.665 391.945 ;
      RECT  138.245 391.585 142.905 391.945 ;
      RECT  144.485 391.585 149.145 391.945 ;
      RECT  150.725 391.585 155.385 391.945 ;
      RECT  156.965 391.585 161.625 391.945 ;
      RECT  163.205 391.585 167.865 391.945 ;
      RECT  169.445 391.585 174.105 391.945 ;
      RECT  175.685 391.585 180.345 391.945 ;
      RECT  181.925 391.585 186.585 391.945 ;
      RECT  188.165 391.585 192.825 391.945 ;
      RECT  194.405 391.585 199.065 391.945 ;
      RECT  200.645 391.585 205.305 391.945 ;
      RECT  206.885 391.585 211.545 391.945 ;
      RECT  213.125 391.585 217.785 391.945 ;
      RECT  219.365 391.585 224.025 391.945 ;
      RECT  225.605 391.585 230.265 391.945 ;
      RECT  231.845 391.585 236.505 391.945 ;
      RECT  238.085 391.585 242.745 391.945 ;
      RECT  244.325 391.585 248.985 391.945 ;
      RECT  250.565 391.585 255.225 391.945 ;
      RECT  256.805 391.585 321.34 391.945 ;
      RECT  341.98 0.62 395.68 0.98 ;
      RECT  368.36 391.585 395.68 391.945 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  322.92 0.98 392.2 2.88 ;
      RECT  322.92 2.88 392.2 389.685 ;
      RECT  322.92 389.685 392.2 391.585 ;
      RECT  392.2 0.98 395.14 2.88 ;
      RECT  392.2 389.685 395.14 391.585 ;
      RECT  395.14 0.98 395.68 2.88 ;
      RECT  395.14 2.88 395.68 389.685 ;
      RECT  395.14 389.685 395.68 391.585 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 389.685 ;
      RECT  2.34 389.685 2.88 391.945 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 389.685 5.82 391.945 ;
      RECT  5.82 0.98 75.94 2.88 ;
      RECT  5.82 2.88 75.94 389.685 ;
      RECT  5.82 389.685 75.94 391.945 ;
   END
END    sky130_sram_1kbytes_1rw1r_20x256_20
END    LIBRARY
