VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_8kbytes_1rw1r_32x2048_32
   CLASS BLOCK ;
   SIZE 1110.54 BY 721.41 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  103.52 0.0 103.9 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  109.36 0.0 109.74 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  115.2 0.0 115.58 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.04 0.0 121.42 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  126.88 0.0 127.26 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.72 0.0 133.1 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  138.56 0.0 138.94 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.4 0.0 144.78 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.24 0.0 150.62 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.08 0.0 156.46 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.92 0.0 162.3 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  167.76 0.0 168.14 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  173.6 0.0 173.98 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.44 0.0 179.82 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  185.28 0.0 185.66 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  191.12 0.0 191.5 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  196.96 0.0 197.34 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  202.8 0.0 203.18 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.64 0.0 209.02 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  214.48 0.0 214.86 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  220.32 0.0 220.7 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.16 0.0 226.54 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.0 0.0 232.38 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  237.84 0.0 238.22 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  243.68 0.0 244.06 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  249.52 0.0 249.9 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.36 0.0 255.74 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.2 0.0 261.58 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.04 0.0 267.42 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  272.88 0.0 273.26 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  278.72 0.0 279.1 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  284.56 0.0 284.94 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  86.0 0.0 86.38 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.84 0.0 92.22 0.38 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.68 0.0 98.06 0.38 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 173.51 0.38 173.89 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 182.01 0.38 182.39 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 187.65 0.38 188.03 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 196.15 0.38 196.53 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 201.79 0.38 202.17 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 210.29 0.38 210.67 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 215.93 0.38 216.31 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 224.43 0.38 224.81 ;
      END
   END addr0[10]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1019.16 721.03 1019.54 721.41 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1013.32 721.03 1013.7 721.41 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1007.48 721.03 1007.86 721.41 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 120.47 1110.54 120.85 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 111.97 1110.54 112.35 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 106.33 1110.54 106.71 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 97.83 1110.54 98.21 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 92.19 1110.54 92.57 ;
      END
   END addr1[7]
   PIN addr1[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 83.69 1110.54 84.07 ;
      END
   END addr1[8]
   PIN addr1[9]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 78.05 1110.54 78.43 ;
      END
   END addr1[9]
   PIN addr1[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  1036.68 0.0 1037.06 0.38 ;
      END
   END addr1[10]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 64.73 0.38 65.11 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 672.385 1110.54 672.765 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 73.23 0.38 73.61 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 65.475 0.38 65.855 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  1110.16 671.695 1110.54 672.075 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  156.77 0.0 157.15 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  181.465 0.0 181.845 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.425 0.0 206.805 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.195 0.0 230.575 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  256.345 0.0 256.725 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  281.305 0.0 281.685 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.265 0.0 306.645 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.225 0.0 331.605 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  356.185 0.0 356.565 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  381.145 0.0 381.525 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  406.105 0.0 406.485 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  431.065 0.0 431.445 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  456.025 0.0 456.405 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  480.985 0.0 481.365 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  505.945 0.0 506.325 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.905 0.0 531.285 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  555.865 0.0 556.245 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  580.825 0.0 581.205 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  605.785 0.0 606.165 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  630.745 0.0 631.125 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  655.705 0.0 656.085 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  680.665 0.0 681.045 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  705.625 0.0 706.005 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  730.585 0.0 730.965 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  755.545 0.0 755.925 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  780.505 0.0 780.885 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  805.465 0.0 805.845 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  830.425 0.0 830.805 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  855.385 0.0 855.765 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  880.345 0.0 880.725 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  905.305 0.0 905.685 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  930.265 0.0 930.645 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  156.565 721.03 156.945 721.41 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  181.525 721.03 181.905 721.41 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.485 721.03 206.865 721.41 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  231.445 721.03 231.825 721.41 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  256.405 721.03 256.785 721.41 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  281.365 721.03 281.745 721.41 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.325 721.03 306.705 721.41 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  331.285 721.03 331.665 721.41 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  356.245 721.03 356.625 721.41 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  381.205 721.03 381.585 721.41 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  406.165 721.03 406.545 721.41 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  431.125 721.03 431.505 721.41 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  456.085 721.03 456.465 721.41 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  481.045 721.03 481.425 721.41 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  506.005 721.03 506.385 721.41 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  530.965 721.03 531.345 721.41 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  555.925 721.03 556.305 721.41 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  580.885 721.03 581.265 721.41 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  605.845 721.03 606.225 721.41 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  630.805 721.03 631.185 721.41 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  655.765 721.03 656.145 721.41 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  680.725 721.03 681.105 721.41 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  705.685 721.03 706.065 721.41 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  730.645 721.03 731.025 721.41 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  755.605 721.03 755.985 721.41 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  780.565 721.03 780.945 721.41 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  805.525 721.03 805.905 721.41 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  830.485 721.03 830.865 721.41 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  855.445 721.03 855.825 721.41 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  880.405 721.03 880.785 721.41 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  905.365 721.03 905.745 721.41 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  930.325 721.03 930.705 721.41 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.74 721.41 ;
         LAYER met4 ;
         RECT  1108.8 0.0 1110.54 721.41 ;
         LAYER met3 ;
         RECT  0.0 0.0 1110.54 1.74 ;
         LAYER met3 ;
         RECT  0.0 719.67 1110.54 721.41 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.48 716.19 1107.06 717.93 ;
         LAYER met3 ;
         RECT  3.48 3.48 1107.06 5.22 ;
         LAYER met4 ;
         RECT  1105.32 3.48 1107.06 717.93 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 717.93 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 1109.92 720.79 ;
   LAYER  met2 ;
      RECT  0.62 0.62 1109.92 720.79 ;
   LAYER  met3 ;
      RECT  0.98 172.91 1109.92 174.49 ;
      RECT  0.62 174.49 0.98 181.41 ;
      RECT  0.62 182.99 0.98 187.05 ;
      RECT  0.62 188.63 0.98 195.55 ;
      RECT  0.62 197.13 0.98 201.19 ;
      RECT  0.62 202.77 0.98 209.69 ;
      RECT  0.62 211.27 0.98 215.33 ;
      RECT  0.62 216.91 0.98 223.83 ;
      RECT  0.98 119.87 1109.56 121.45 ;
      RECT  0.98 121.45 1109.56 172.91 ;
      RECT  1109.56 121.45 1109.92 172.91 ;
      RECT  1109.56 112.95 1109.92 119.87 ;
      RECT  1109.56 107.31 1109.92 111.37 ;
      RECT  1109.56 98.81 1109.92 105.73 ;
      RECT  1109.56 93.17 1109.92 97.23 ;
      RECT  1109.56 84.67 1109.92 91.59 ;
      RECT  1109.56 79.03 1109.92 83.09 ;
      RECT  0.98 174.49 1109.56 671.785 ;
      RECT  0.98 671.785 1109.56 673.365 ;
      RECT  0.62 74.21 0.98 172.91 ;
      RECT  0.62 66.455 0.98 72.63 ;
      RECT  1109.56 174.49 1109.92 671.095 ;
      RECT  1109.56 2.34 1109.92 77.45 ;
      RECT  0.62 2.34 0.98 64.13 ;
      RECT  0.62 225.41 0.98 719.07 ;
      RECT  1109.56 673.365 1109.92 719.07 ;
      RECT  0.98 673.365 2.88 715.59 ;
      RECT  0.98 715.59 2.88 718.53 ;
      RECT  0.98 718.53 2.88 719.07 ;
      RECT  2.88 673.365 1107.66 715.59 ;
      RECT  2.88 718.53 1107.66 719.07 ;
      RECT  1107.66 673.365 1109.56 715.59 ;
      RECT  1107.66 715.59 1109.56 718.53 ;
      RECT  1107.66 718.53 1109.56 719.07 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 119.87 ;
      RECT  2.88 2.34 1107.66 2.88 ;
      RECT  2.88 5.82 1107.66 119.87 ;
      RECT  1107.66 2.34 1109.56 2.88 ;
      RECT  1107.66 2.88 1109.56 5.82 ;
      RECT  1107.66 5.82 1109.56 119.87 ;
   LAYER  met4 ;
      RECT  102.92 0.98 104.5 720.79 ;
      RECT  104.5 0.62 108.76 0.98 ;
      RECT  110.34 0.62 114.6 0.98 ;
      RECT  116.18 0.62 120.44 0.98 ;
      RECT  122.02 0.62 126.28 0.98 ;
      RECT  127.86 0.62 132.12 0.98 ;
      RECT  133.7 0.62 137.96 0.98 ;
      RECT  139.54 0.62 143.8 0.98 ;
      RECT  145.38 0.62 149.64 0.98 ;
      RECT  151.22 0.62 155.48 0.98 ;
      RECT  162.9 0.62 167.16 0.98 ;
      RECT  168.74 0.62 173.0 0.98 ;
      RECT  174.58 0.62 178.84 0.98 ;
      RECT  186.26 0.62 190.52 0.98 ;
      RECT  192.1 0.62 196.36 0.98 ;
      RECT  197.94 0.62 202.2 0.98 ;
      RECT  209.62 0.62 213.88 0.98 ;
      RECT  215.46 0.62 219.72 0.98 ;
      RECT  221.3 0.62 225.56 0.98 ;
      RECT  232.98 0.62 237.24 0.98 ;
      RECT  238.82 0.62 243.08 0.98 ;
      RECT  244.66 0.62 248.92 0.98 ;
      RECT  250.5 0.62 254.76 0.98 ;
      RECT  262.18 0.62 266.44 0.98 ;
      RECT  268.02 0.62 272.28 0.98 ;
      RECT  273.86 0.62 278.12 0.98 ;
      RECT  86.98 0.62 91.24 0.98 ;
      RECT  92.82 0.62 97.08 0.98 ;
      RECT  98.66 0.62 102.92 0.98 ;
      RECT  104.5 0.98 1018.56 720.43 ;
      RECT  1018.56 0.98 1020.14 720.43 ;
      RECT  1014.3 720.43 1018.56 720.79 ;
      RECT  1008.46 720.43 1012.72 720.79 ;
      RECT  157.75 0.62 161.32 0.98 ;
      RECT  180.42 0.62 180.865 0.98 ;
      RECT  182.445 0.62 184.68 0.98 ;
      RECT  203.78 0.62 205.825 0.98 ;
      RECT  207.405 0.62 208.04 0.98 ;
      RECT  227.14 0.62 229.595 0.98 ;
      RECT  231.175 0.62 231.4 0.98 ;
      RECT  257.325 0.62 260.6 0.98 ;
      RECT  279.7 0.62 280.705 0.98 ;
      RECT  282.285 0.62 283.96 0.98 ;
      RECT  285.54 0.62 305.665 0.98 ;
      RECT  307.245 0.62 330.625 0.98 ;
      RECT  332.205 0.62 355.585 0.98 ;
      RECT  357.165 0.62 380.545 0.98 ;
      RECT  382.125 0.62 405.505 0.98 ;
      RECT  407.085 0.62 430.465 0.98 ;
      RECT  432.045 0.62 455.425 0.98 ;
      RECT  457.005 0.62 480.385 0.98 ;
      RECT  481.965 0.62 505.345 0.98 ;
      RECT  506.925 0.62 530.305 0.98 ;
      RECT  531.885 0.62 555.265 0.98 ;
      RECT  556.845 0.62 580.225 0.98 ;
      RECT  581.805 0.62 605.185 0.98 ;
      RECT  606.765 0.62 630.145 0.98 ;
      RECT  631.725 0.62 655.105 0.98 ;
      RECT  656.685 0.62 680.065 0.98 ;
      RECT  681.645 0.62 705.025 0.98 ;
      RECT  706.605 0.62 729.985 0.98 ;
      RECT  731.565 0.62 754.945 0.98 ;
      RECT  756.525 0.62 779.905 0.98 ;
      RECT  781.485 0.62 804.865 0.98 ;
      RECT  806.445 0.62 829.825 0.98 ;
      RECT  831.405 0.62 854.785 0.98 ;
      RECT  856.365 0.62 879.745 0.98 ;
      RECT  881.325 0.62 904.705 0.98 ;
      RECT  906.285 0.62 929.665 0.98 ;
      RECT  931.245 0.62 1036.08 0.98 ;
      RECT  104.5 720.43 155.965 720.79 ;
      RECT  157.545 720.43 180.925 720.79 ;
      RECT  182.505 720.43 205.885 720.79 ;
      RECT  207.465 720.43 230.845 720.79 ;
      RECT  232.425 720.43 255.805 720.79 ;
      RECT  257.385 720.43 280.765 720.79 ;
      RECT  282.345 720.43 305.725 720.79 ;
      RECT  307.305 720.43 330.685 720.79 ;
      RECT  332.265 720.43 355.645 720.79 ;
      RECT  357.225 720.43 380.605 720.79 ;
      RECT  382.185 720.43 405.565 720.79 ;
      RECT  407.145 720.43 430.525 720.79 ;
      RECT  432.105 720.43 455.485 720.79 ;
      RECT  457.065 720.43 480.445 720.79 ;
      RECT  482.025 720.43 505.405 720.79 ;
      RECT  506.985 720.43 530.365 720.79 ;
      RECT  531.945 720.43 555.325 720.79 ;
      RECT  556.905 720.43 580.285 720.79 ;
      RECT  581.865 720.43 605.245 720.79 ;
      RECT  606.825 720.43 630.205 720.79 ;
      RECT  631.785 720.43 655.165 720.79 ;
      RECT  656.745 720.43 680.125 720.79 ;
      RECT  681.705 720.43 705.085 720.79 ;
      RECT  706.665 720.43 730.045 720.79 ;
      RECT  731.625 720.43 755.005 720.79 ;
      RECT  756.585 720.43 779.965 720.79 ;
      RECT  781.545 720.43 804.925 720.79 ;
      RECT  806.505 720.43 829.885 720.79 ;
      RECT  831.465 720.43 854.845 720.79 ;
      RECT  856.425 720.43 879.805 720.79 ;
      RECT  881.385 720.43 904.765 720.79 ;
      RECT  906.345 720.43 929.725 720.79 ;
      RECT  931.305 720.43 1006.88 720.79 ;
      RECT  2.34 0.62 85.4 0.98 ;
      RECT  1020.14 720.43 1108.2 720.79 ;
      RECT  1037.66 0.62 1108.2 0.98 ;
      RECT  1020.14 0.98 1104.72 2.88 ;
      RECT  1020.14 2.88 1104.72 718.53 ;
      RECT  1020.14 718.53 1104.72 720.43 ;
      RECT  1104.72 0.98 1107.66 2.88 ;
      RECT  1104.72 718.53 1107.66 720.43 ;
      RECT  1107.66 0.98 1108.2 2.88 ;
      RECT  1107.66 2.88 1108.2 718.53 ;
      RECT  1107.66 718.53 1108.2 720.43 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 718.53 ;
      RECT  2.34 718.53 2.88 720.79 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 718.53 5.82 720.79 ;
      RECT  5.82 0.98 102.92 2.88 ;
      RECT  5.82 2.88 102.92 718.53 ;
      RECT  5.82 718.53 102.92 720.79 ;
   END
END    sky130_sram_8kbytes_1rw1r_32x2048_32
END    LIBRARY
